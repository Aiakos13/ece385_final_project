module sprite_table(input logic frame_clk,
						  input logic [7:0] last_key_code,
						  input logic [9:0] X, Y,
						 // input int hunger,happiness,
						  output logic [31:0] color);
/*						  
#include <stdint.h>

#define MAIN_CHARACTER JODI_FRAME_COUNT 4
#define MAIN_CHARACTER JODI_FRAME_WIDTH 100
#define MAIN_CHARACTER JODI_FRAME_HEIGHT 100

// Piskel data for "Main Character Jodi" 

static const uint32_t main_character jodi_data[4][10000] = {
{*/
logic [9:0] Xval,Yval;//,B1X,B1Y,B2X,B2Y;


logic [31:0] jodi_left[1024];
logic [31:0] jodi_right[1024];
logic [31:0] jodi_up[1024];
logic [31:0] jodi_down[1024];
/*
logic [7:0] last_key_code;

always_ff @(posedge frame_clk)
begin
	if (sprite == 8'h50 || sprite == 8'h4F || sprite == 8'h52 || sprite == 8'h51)
		last_key_code <= sprite;
	else
		last_key_code <= last_key_code;
end
*/
always_comb
begin
jodi_left = '{
32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 
32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 
32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 
32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 
32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'hff191919, 32'hff191919, 32'h00000000, 32'h00000000, 32'h00000000, 32'hff191919, 32'hff191919, 32'hff191919, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 
32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'hff191919, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'hff191919, 32'hffb002d7, 32'hffb002d7, 32'hff191919, 32'h00000000, 32'hff191919, 32'hffb002d7, 32'hffb002d7, 32'hffb002d7, 32'hff191919, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 
32'h00000000, 32'h00000000, 32'h00000000, 32'hff191919, 32'hff191919, 32'hff191919, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'hff191919, 32'hffb002d7, 32'hffb002d7, 32'hffb002d7, 32'hff191919, 32'hff191919, 32'hffb002d7, 32'hffb002d7, 32'hffb002d7, 32'hffb002d7, 32'hff191919, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 
32'h00000000, 32'h00000000, 32'h00000000, 32'hff191919, 32'hffb002d7, 32'hff191919, 32'hff191919, 32'hff191919, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'hff191919, 32'hffb002d7, 32'hffb002d7, 32'hffb002d7, 32'hffb002d7, 32'hffb002d7, 32'hffb002d7, 32'hff191919, 32'hff191919, 32'hff191919, 32'hff191919, 32'hff191919, 32'hff191919, 32'hff191919, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 
32'h00000000, 32'h00000000, 32'h00000000, 32'hff191919, 32'hffb002d7, 32'hffb002d7, 32'hffd8dc29, 32'hff191919, 32'h00000000, 32'h00000000, 32'hff191919, 32'hff191919, 32'hff191919, 32'hff191919, 32'hffb002d7, 32'hffb002d7, 32'hffb002d7, 32'hffb002d7, 32'hffb002d7, 32'hffb002d7, 32'hff191919, 32'hffd8dc29, 32'hffd8dc29, 32'hffd8dc29, 32'hffd8dc29, 32'hff191919, 32'hff191919, 32'hff191919, 32'hff191919, 32'h00000000, 32'h00000000, 32'h00000000, 
32'h00000000, 32'h00000000, 32'h00000000, 32'hff191919, 32'hffd8dc29, 32'hffd8dc29, 32'hffb002d7, 32'hff191919, 32'h00000000, 32'hff191919, 32'hff191919, 32'hffd8dc29, 32'hffd8dc29, 32'hff191919, 32'hffb002d7, 32'hffb002d7, 32'hffb002d7, 32'hffb002d7, 32'hffb002d7, 32'hffb002d7, 32'hff191919, 32'hffd8dc29, 32'hffd8dc29, 32'hffd8dc29, 32'hff191919, 32'hffd8dc29, 32'hffd8dc29, 32'hffd8dc29, 32'hffd8dc29, 32'hff191919, 32'h00000000, 32'h00000000, 
32'h00000000, 32'h00000000, 32'h00000000, 32'hff191919, 32'hffb002d7, 32'hffd8dc29, 32'hffd8dc29, 32'hffd8dc29, 32'hff191919, 32'hff191919, 32'hffd8dc29, 32'hffd8dc29, 32'hffd8dc29, 32'hff191919, 32'hffb002d7, 32'hffb002d7, 32'hffb002d7, 32'hffb002d7, 32'hffb002d7, 32'hffb002d7, 32'hffb002d7, 32'hff191919, 32'hffd8dc29, 32'hff191919, 32'hffd8dc29, 32'hffd8dc29, 32'hffd8dc29, 32'hffd8dc29, 32'hffd8dc29, 32'hffd8dc29, 32'hff191919, 32'h00000000, 
32'h00000000, 32'h00000000, 32'h00000000, 32'hff191919, 32'hffd8dc29, 32'hffb002d7, 32'hffb002d7, 32'hffb002d7, 32'hffb002d7, 32'hffd8dc29, 32'hffd8dc29, 32'hffd8dc29, 32'hffd8dc29, 32'hffd8dc29, 32'hff191919, 32'hffb002d7, 32'hffb002d7, 32'hffb002d7, 32'hffb002d7, 32'hffb002d7, 32'hffb002d7, 32'hffd8dc29, 32'hffd8dc29, 32'hffd8dc29, 32'hffd8dc29, 32'hffd8dc29, 32'hffd8dc29, 32'hffd8dc29, 32'hffd8dc29, 32'hffd8dc29, 32'hff191919, 32'h00000000, 
32'h00000000, 32'h00000000, 32'h00000000, 32'hff191919, 32'hffd8dc29, 32'hffd8dc29, 32'hffd8dc29, 32'hffd8dc29, 32'hffd8dc29, 32'hffd8dc29, 32'hffd8dc29, 32'hffd8dc29, 32'hffd8dc29, 32'hffd8dc29, 32'hffd8dc29, 32'hff191919, 32'hff191919, 32'hffb002d7, 32'hffb002d7, 32'hffb002d7, 32'hffd8dc29, 32'hffd8dc29, 32'hffd8dc29, 32'hff191919, 32'hff191919, 32'hff191919, 32'hffd8dc29, 32'hffd8dc29, 32'hff191919, 32'hff191919, 32'h00000000, 32'h00000000, 
32'h00000000, 32'h00000000, 32'h00000000, 32'hff191919, 32'hffd8dc29, 32'hffb002d7, 32'hffb002d7, 32'hffb002d7, 32'hffb002d7, 32'hffd8dc29, 32'hffd8dc29, 32'hffd8dc29, 32'hffd8dc29, 32'hffd8dc29, 32'hffd8dc29, 32'hffd8dc29, 32'hff191919, 32'hffb002d7, 32'hffb002d7, 32'hffd8dc29, 32'hffd8dc29, 32'hffd8dc29, 32'hff191919, 32'hffffffff, 32'hff191919, 32'hff191919, 32'hffd8dc29, 32'hffd8dc29, 32'hff191919, 32'h00000000, 32'h00000000, 32'h00000000, 
32'h00000000, 32'h00000000, 32'h00000000, 32'hff191919, 32'hffd8dc29, 32'hffb002d7, 32'hffd8dc29, 32'hffd8dc29, 32'hffd8dc29, 32'hffd8dc29, 32'hffd8dc29, 32'hffd8dc29, 32'hffd8dc29, 32'hffd8dc29, 32'hffd8dc29, 32'hffd8dc29, 32'hff191919, 32'hff191919, 32'hffd8dc29, 32'hffd8dc29, 32'hffd8dc29, 32'hffd8dc29, 32'hff191919, 32'hffffffff, 32'hff191919, 32'hff191919, 32'hffd8dc29, 32'hffd8dc29, 32'hff191919, 32'h00000000, 32'h00000000, 32'h00000000, 
32'h00000000, 32'h00000000, 32'h00000000, 32'hff191919, 32'hffb002d7, 32'hffb002d7, 32'hffd8dc29, 32'hffb002d7, 32'hffb002d7, 32'hffd8dc29, 32'hffd8dc29, 32'hffd8dc29, 32'hffd8dc29, 32'hffd8dc29, 32'hffd8dc29, 32'hffd8dc29, 32'hffd8dc29, 32'hffd8dc29, 32'hffd8dc29, 32'hffd8dc29, 32'hffd8dc29, 32'hffd8dc29, 32'hff191919, 32'hffffffff, 32'hffffffff, 32'hff191919, 32'hffd8dc29, 32'hffd8dc29, 32'hff191919, 32'h00000000, 32'h00000000, 32'h00000000, 
32'h00000000, 32'h00000000, 32'h00000000, 32'hff191919, 32'hffd8dc29, 32'hffd8dc29, 32'hffd8dc29, 32'hffb002d7, 32'hff191919, 32'hff191919, 32'hffd8dc29, 32'hffd8dc29, 32'hffd8dc29, 32'hffd8dc29, 32'hffd8dc29, 32'hffd8dc29, 32'hffd8dc29, 32'hffd8dc29, 32'hffd8dc29, 32'hffd8dc29, 32'hffd8dc29, 32'hffd8dc29, 32'hffd8dc29, 32'hff191919, 32'hff191919, 32'hff191919, 32'hffd8dc29, 32'hff191919, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 
32'h00000000, 32'h00000000, 32'h00000000, 32'hff191919, 32'hffd8dc29, 32'hffd8dc29, 32'hffb002d7, 32'hffb002d7, 32'hff191919, 32'h00000000, 32'hff191919, 32'hffd8dc29, 32'hffd8dc29, 32'hffd8dc29, 32'hffd8dc29, 32'hffd8dc29, 32'hffd8dc29, 32'hffd8dc29, 32'hffd8dc29, 32'hffd8dc29, 32'hffd8dc29, 32'hffd8dc29, 32'hffd8dc29, 32'hffd8dc29, 32'hffd8dc29, 32'hffd8dc29, 32'hff191919, 32'hff191919, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 
32'h00000000, 32'h00000000, 32'h00000000, 32'hff191919, 32'hffb002d7, 32'hffb002d7, 32'hffb002d7, 32'hff191919, 32'h00000000, 32'h00000000, 32'h00000000, 32'hff191919, 32'hffd8dc29, 32'hffd8dc29, 32'hffd8dc29, 32'hffd8dc29, 32'hffb002d7, 32'hffb002d7, 32'hffb002d7, 32'hffb002d7, 32'hffd8dc29, 32'hffd8dc29, 32'hffd8dc29, 32'hffd8dc29, 32'hff191919, 32'hff191919, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 
32'h00000000, 32'h00000000, 32'h00000000, 32'hff191919, 32'hffb002d7, 32'hff191919, 32'hff191919, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'hff191919, 32'hff191919, 32'hff191919, 32'hffd8dc29, 32'hffb002d7, 32'hffb002d7, 32'hffb002d7, 32'hffb002d7, 32'hffb002d7, 32'hffb002d7, 32'hffd8dc29, 32'hff191919, 32'hff191919, 32'hff191919, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 
32'h00000000, 32'h00000000, 32'h00000000, 32'hff191919, 32'hff191919, 32'hff191919, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'hff191919, 32'hff191919, 32'hffb002d7, 32'hffb002d7, 32'hffb002d7, 32'hffb002d7, 32'hffb002d7, 32'hffb002d7, 32'hff191919, 32'hff191919, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 
32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'hff191919, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'hff191919, 32'hffb002d7, 32'hffb002d7, 32'hffb002d7, 32'hffb002d7, 32'hffb002d7, 32'hffb002d7, 32'hff191919, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 
32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'hff191919, 32'hffb002d7, 32'hffb002d7, 32'hffb002d7, 32'hffb002d7, 32'hffb002d7, 32'hff191919, 32'hff191919, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 
32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'hff191919, 32'hffb002d7, 32'hffb002d7, 32'hffb002d7, 32'hffb002d7, 32'hff191919, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 
32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'hff191919, 32'hffb002d7, 32'hffb002d7, 32'hffb002d7, 32'hffb002d7, 32'hff191919, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 
32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'hff191919, 32'hff191919, 32'hff191919, 32'hff191919, 32'hff191919, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 
32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 
32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 
32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 
32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 
32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 
32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000
};
jodi_right = '{
32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 
32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 
32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 
32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 
32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 
32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 
32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'hff191919, 32'hff191919, 32'hff191919, 32'h00000000, 32'h00000000, 32'h00000000, 32'hff191919, 32'hff191919, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 
32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'hff191919, 32'hffb002d7, 32'hffb002d7, 32'hffb002d7, 32'hff191919, 32'h00000000, 32'hff191919, 32'hffb002d7, 32'hffb002d7, 32'hff191919, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'hff191919, 32'h00000000, 32'h00000000, 32'h00000000, 
32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'hff191919, 32'hffb002d7, 32'hffb002d7, 32'hffb002d7, 32'hffb002d7, 32'hff191919, 32'hff191919, 32'hffb002d7, 32'hffb002d7, 32'hffb002d7, 32'hff191919, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'hff191919, 32'hff191919, 32'hff191919, 32'h00000000, 32'h00000000, 
32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'hff191919, 32'hff191919, 32'hff191919, 32'hff191919, 32'hff191919, 32'hff191919, 32'hff191919, 32'hffb002d7, 32'hffb002d7, 32'hffb002d7, 32'hffb002d7, 32'hffb002d7, 32'hffb002d7, 32'hff191919, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'hff191919, 32'hff191919, 32'hff191919, 32'hffb002d7, 32'hff191919, 32'h00000000, 32'h00000000, 
32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'hff191919, 32'hff191919, 32'hff191919, 32'hff191919, 32'hffd8dc29, 32'hffd8dc29, 32'hffd8dc29, 32'hffd8dc29, 32'hff191919, 32'hffb002d7, 32'hffb002d7, 32'hffb002d7, 32'hffb002d7, 32'hffb002d7, 32'hffb002d7, 32'hff191919, 32'hff191919, 32'hff191919, 32'hff191919, 32'h00000000, 32'h00000000, 32'hff191919, 32'hffd8dc29, 32'hffb002d7, 32'hffb002d7, 32'hff191919, 32'h00000000, 32'h00000000, 
32'h00000000, 32'h00000000, 32'h00000000, 32'hff191919, 32'hffd8dc29, 32'hffd8dc29, 32'hffd8dc29, 32'hffd8dc29, 32'hff191919, 32'hffd8dc29, 32'hffd8dc29, 32'hffd8dc29, 32'hff191919, 32'hffb002d7, 32'hffb002d7, 32'hffb002d7, 32'hffb002d7, 32'hffb002d7, 32'hffb002d7, 32'hff191919, 32'hffd8dc29, 32'hffd8dc29, 32'hff191919, 32'hff191919, 32'h00000000, 32'hff191919, 32'hffb002d7, 32'hffd8dc29, 32'hffd8dc29, 32'hff191919, 32'h00000000, 32'h00000000, 
32'h00000000, 32'h00000000, 32'hff191919, 32'hffd8dc29, 32'hffd8dc29, 32'hffd8dc29, 32'hffd8dc29, 32'hffd8dc29, 32'hffd8dc29, 32'hff191919, 32'hffd8dc29, 32'hff191919, 32'hffb002d7, 32'hffb002d7, 32'hffb002d7, 32'hffb002d7, 32'hffb002d7, 32'hffb002d7, 32'hffb002d7, 32'hff191919, 32'hffd8dc29, 32'hffd8dc29, 32'hffd8dc29, 32'hff191919, 32'hff191919, 32'hffd8dc29, 32'hffd8dc29, 32'hffd8dc29, 32'hffb002d7, 32'hff191919, 32'h00000000, 32'h00000000, 
32'h00000000, 32'h00000000, 32'hff191919, 32'hffd8dc29, 32'hffd8dc29, 32'hffd8dc29, 32'hffd8dc29, 32'hffd8dc29, 32'hffd8dc29, 32'hffd8dc29, 32'hffd8dc29, 32'hffd8dc29, 32'hffb002d7, 32'hffb002d7, 32'hffb002d7, 32'hffb002d7, 32'hffb002d7, 32'hffb002d7, 32'hff191919, 32'hffd8dc29, 32'hffd8dc29, 32'hffd8dc29, 32'hffd8dc29, 32'hffd8dc29, 32'hffb002d7, 32'hffb002d7, 32'hffb002d7, 32'hffb002d7, 32'hffd8dc29, 32'hff191919, 32'h00000000, 32'h00000000, 
32'h00000000, 32'h00000000, 32'h00000000, 32'hff191919, 32'hff191919, 32'hffd8dc29, 32'hffd8dc29, 32'hff191919, 32'hff191919, 32'hff191919, 32'hffd8dc29, 32'hffd8dc29, 32'hffd8dc29, 32'hffb002d7, 32'hffb002d7, 32'hffb002d7, 32'hff191919, 32'hff191919, 32'hffd8dc29, 32'hffd8dc29, 32'hffd8dc29, 32'hffd8dc29, 32'hffd8dc29, 32'hffd8dc29, 32'hffd8dc29, 32'hffd8dc29, 32'hffd8dc29, 32'hffd8dc29, 32'hffd8dc29, 32'hff191919, 32'h00000000, 32'h00000000, 
32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'hff191919, 32'hffd8dc29, 32'hffd8dc29, 32'hff191919, 32'hff191919, 32'hffffffff, 32'hff191919, 32'hffd8dc29, 32'hffd8dc29, 32'hffd8dc29, 32'hffb002d7, 32'hffb002d7, 32'hff191919, 32'hffd8dc29, 32'hffd8dc29, 32'hffd8dc29, 32'hffd8dc29, 32'hffd8dc29, 32'hffd8dc29, 32'hffd8dc29, 32'hffb002d7, 32'hffb002d7, 32'hffb002d7, 32'hffb002d7, 32'hffd8dc29, 32'hff191919, 32'h00000000, 32'h00000000, 
32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'hff191919, 32'hffd8dc29, 32'hffd8dc29, 32'hff191919, 32'hff191919, 32'hffffffff, 32'hff191919, 32'hffd8dc29, 32'hffd8dc29, 32'hffd8dc29, 32'hffd8dc29, 32'hff191919, 32'hff191919, 32'hffd8dc29, 32'hffd8dc29, 32'hffd8dc29, 32'hffd8dc29, 32'hffd8dc29, 32'hffd8dc29, 32'hffd8dc29, 32'hffd8dc29, 32'hffd8dc29, 32'hffd8dc29, 32'hffb002d7, 32'hffd8dc29, 32'hff191919, 32'h00000000, 32'h00000000, 
32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'hff191919, 32'hffd8dc29, 32'hffd8dc29, 32'hff191919, 32'hffffffff, 32'hffffffff, 32'hff191919, 32'hffd8dc29, 32'hffd8dc29, 32'hffd8dc29, 32'hffd8dc29, 32'hffd8dc29, 32'hffd8dc29, 32'hffd8dc29, 32'hffd8dc29, 32'hffd8dc29, 32'hffd8dc29, 32'hffd8dc29, 32'hffd8dc29, 32'hffd8dc29, 32'hffb002d7, 32'hffb002d7, 32'hffd8dc29, 32'hffb002d7, 32'hffb002d7, 32'hff191919, 32'h00000000, 32'h00000000, 
32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'hff191919, 32'hffd8dc29, 32'hff191919, 32'hff191919, 32'hff191919, 32'hffd8dc29, 32'hffd8dc29, 32'hffd8dc29, 32'hffd8dc29, 32'hffd8dc29, 32'hffd8dc29, 32'hffd8dc29, 32'hffd8dc29, 32'hffd8dc29, 32'hffd8dc29, 32'hffd8dc29, 32'hffd8dc29, 32'hffd8dc29, 32'hff191919, 32'hff191919, 32'hffb002d7, 32'hffd8dc29, 32'hffd8dc29, 32'hffd8dc29, 32'hff191919, 32'h00000000, 32'h00000000, 
32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'hff191919, 32'hff191919, 32'hffd8dc29, 32'hffd8dc29, 32'hffd8dc29, 32'hffd8dc29, 32'hffd8dc29, 32'hffd8dc29, 32'hffd8dc29, 32'hffd8dc29, 32'hffd8dc29, 32'hffd8dc29, 32'hffd8dc29, 32'hffd8dc29, 32'hffd8dc29, 32'hffd8dc29, 32'hffd8dc29, 32'hff191919, 32'h00000000, 32'hff191919, 32'hffb002d7, 32'hffb002d7, 32'hffd8dc29, 32'hffd8dc29, 32'hff191919, 32'h00000000, 32'h00000000, 
32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'hff191919, 32'hff191919, 32'hffd8dc29, 32'hffd8dc29, 32'hffd8dc29, 32'hffd8dc29, 32'hffb002d7, 32'hffb002d7, 32'hffb002d7, 32'hffb002d7, 32'hffd8dc29, 32'hffd8dc29, 32'hffd8dc29, 32'hffd8dc29, 32'hff191919, 32'h00000000, 32'h00000000, 32'h00000000, 32'hff191919, 32'hffb002d7, 32'hffb002d7, 32'hffb002d7, 32'hff191919, 32'h00000000, 32'h00000000, 
32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'hff191919, 32'hff191919, 32'hff191919, 32'hffd8dc29, 32'hffb002d7, 32'hffb002d7, 32'hffb002d7, 32'hffb002d7, 32'hffb002d7, 32'hffb002d7, 32'hffd8dc29, 32'hff191919, 32'hff191919, 32'hff191919, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'hff191919, 32'hff191919, 32'hffb002d7, 32'hff191919, 32'h00000000, 32'h00000000, 
32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'hff191919, 32'hff191919, 32'hffb002d7, 32'hffb002d7, 32'hffb002d7, 32'hffb002d7, 32'hffb002d7, 32'hffb002d7, 32'hff191919, 32'hff191919, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'hff191919, 32'hff191919, 32'hff191919, 32'h00000000, 32'h00000000, 
32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'hff191919, 32'hffb002d7, 32'hffb002d7, 32'hffb002d7, 32'hffb002d7, 32'hffb002d7, 32'hffb002d7, 32'hff191919, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'hff191919, 32'h00000000, 32'h00000000, 32'h00000000, 
32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'hff191919, 32'hff191919, 32'hffb002d7, 32'hffb002d7, 32'hffb002d7, 32'hffb002d7, 32'hffb002d7, 32'hff191919, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 
32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'hff191919, 32'hffb002d7, 32'hffb002d7, 32'hffb002d7, 32'hffb002d7, 32'hff191919, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 
32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'hff191919, 32'hffb002d7, 32'hffb002d7, 32'hffb002d7, 32'hffb002d7, 32'hff191919, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 
32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'hff191919, 32'hff191919, 32'hff191919, 32'hff191919, 32'hff191919, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 
32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 
32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 
32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 
32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000
};
jodi_up = '{
32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'hff191919, 32'hff191919, 32'hff191919, 32'hff191919, 32'hff191919, 32'hff191919, 32'hff191919, 32'hff191919, 32'hff191919, 32'hff191919, 32'hff191919, 32'hff191919, 32'hff191919, 32'hff191919, 32'hff191919, 32'hff191919, 32'hff191919, 32'hff191919, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 
32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'hff191919, 32'hff191919, 32'hffb002d7, 32'hffb002d7, 32'hffd8dc29, 32'hffd8dc29, 32'hffd8dc29, 32'hffb002d7, 32'hffb002d7, 32'hffd8dc29, 32'hffb002d7, 32'hffb002d7, 32'hffd8dc29, 32'hffb002d7, 32'hffb002d7, 32'hffb002d7, 32'hff191919, 32'hff191919, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 
32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'hff191919, 32'hff191919, 32'hffb002d7, 32'hffb002d7, 32'hffd8dc29, 32'hffb002d7, 32'hffb002d7, 32'hffd8dc29, 32'hffb002d7, 32'hffb002d7, 32'hffd8dc29, 32'hffb002d7, 32'hff191919, 32'hff191919, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 
32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'hff191919, 32'hff191919, 32'hffd8dc29, 32'hffd8dc29, 32'hffb002d7, 32'hffd8dc29, 32'hffb002d7, 32'hffd8dc29, 32'hff191919, 32'hff191919, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 
32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'hff191919, 32'hff191919, 32'hff191919, 32'hffd8dc29, 32'hffd8dc29, 32'hff191919, 32'hff191919, 32'hff191919, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 
32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'hff191919, 32'hffd8dc29, 32'hffd8dc29, 32'hff191919, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 
32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'hff191919, 32'hff191919, 32'hffd8dc29, 32'hffd8dc29, 32'hff191919, 32'hff191919, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 
32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'hff191919, 32'hff191919, 32'hffd8dc29, 32'hffd8dc29, 32'hffd8dc29, 32'hffd8dc29, 32'hff191919, 32'hff191919, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 
32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'hff191919, 32'hff191919, 32'hffd8dc29, 32'hffd8dc29, 32'hffd8dc29, 32'hffd8dc29, 32'hffd8dc29, 32'hffd8dc29, 32'hff191919, 32'hff191919, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 
32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'hff191919, 32'hff191919, 32'hffd8dc29, 32'hffd8dc29, 32'hffd8dc29, 32'hff191919, 32'hff191919, 32'hffd8dc29, 32'hffd8dc29, 32'hffd8dc29, 32'hff191919, 32'hff191919, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 
32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'hff191919, 32'hff191919, 32'hffd8dc29, 32'hffd8dc29, 32'hffd8dc29, 32'hff191919, 32'hff191919, 32'hff191919, 32'hff191919, 32'hffd8dc29, 32'hffd8dc29, 32'hffd8dc29, 32'hff191919, 32'hff191919, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 
32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'hff191919, 32'hff191919, 32'hff191919, 32'hff191919, 32'hffd8dc29, 32'hffd8dc29, 32'hffd8dc29, 32'hffd8dc29, 32'hff191919, 32'hffb002d7, 32'hffb002d7, 32'hff191919, 32'hffd8dc29, 32'hffd8dc29, 32'hffd8dc29, 32'hffd8dc29, 32'hff191919, 32'hff191919, 32'hff191919, 32'hff191919, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 
32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'hff191919, 32'hff191919, 32'hff191919, 32'hffb002d7, 32'hff191919, 32'hffd8dc29, 32'hffd8dc29, 32'hffd8dc29, 32'hffd8dc29, 32'hffd8dc29, 32'hff191919, 32'hffb002d7, 32'hffb002d7, 32'hff191919, 32'hffd8dc29, 32'hffd8dc29, 32'hffd8dc29, 32'hffd8dc29, 32'hffd8dc29, 32'hff191919, 32'hffb002d7, 32'hff191919, 32'hff191919, 32'hff191919, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 
32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'hff191919, 32'hffb002d7, 32'hffb002d7, 32'hffb002d7, 32'hff191919, 32'hffd8dc29, 32'hffd8dc29, 32'hffd8dc29, 32'hffd8dc29, 32'hff191919, 32'hff191919, 32'hffb002d7, 32'hffb002d7, 32'hff191919, 32'hff191919, 32'hffd8dc29, 32'hffd8dc29, 32'hffd8dc29, 32'hffd8dc29, 32'hff191919, 32'hffb002d7, 32'hffb002d7, 32'hffb002d7, 32'hff191919, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 
32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'hff191919, 32'hffb002d7, 32'hffb002d7, 32'hffb002d7, 32'hff191919, 32'hffd8dc29, 32'hffd8dc29, 32'hffd8dc29, 32'hffd8dc29, 32'hff191919, 32'hffb002d7, 32'hffb002d7, 32'hffb002d7, 32'hffb002d7, 32'hff191919, 32'hffd8dc29, 32'hffd8dc29, 32'hffd8dc29, 32'hffd8dc29, 32'hff191919, 32'hffb002d7, 32'hffb002d7, 32'hffb002d7, 32'hff191919, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 
32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'hff191919, 32'hff191919, 32'hffb002d7, 32'hffb002d7, 32'hff191919, 32'hffd8dc29, 32'hffd8dc29, 32'hffd8dc29, 32'hffd8dc29, 32'hff191919, 32'hffb002d7, 32'hffb002d7, 32'hffb002d7, 32'hffb002d7, 32'hff191919, 32'hffd8dc29, 32'hffd8dc29, 32'hffd8dc29, 32'hffd8dc29, 32'hff191919, 32'hffb002d7, 32'hffb002d7, 32'hff191919, 32'hff191919, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 
32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'hff191919, 32'hffb002d7, 32'hffb002d7, 32'hff191919, 32'hffd8dc29, 32'hffd8dc29, 32'hffd8dc29, 32'hffd8dc29, 32'hff191919, 32'hffb002d7, 32'hffb002d7, 32'hffb002d7, 32'hffb002d7, 32'hff191919, 32'hffd8dc29, 32'hffd8dc29, 32'hffd8dc29, 32'hffd8dc29, 32'hff191919, 32'hffb002d7, 32'hffb002d7, 32'hff191919, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 
32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'hff191919, 32'hffb002d7, 32'hffb002d7, 32'hff191919, 32'hffd8dc29, 32'hffd8dc29, 32'hffd8dc29, 32'hffd8dc29, 32'hff191919, 32'hffb002d7, 32'hffb002d7, 32'hffb002d7, 32'hffb002d7, 32'hff191919, 32'hffd8dc29, 32'hffd8dc29, 32'hffd8dc29, 32'hffd8dc29, 32'hff191919, 32'hffb002d7, 32'hffb002d7, 32'hff191919, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 
32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'hff191919, 32'hff191919, 32'hffb002d7, 32'hff191919, 32'hffd8dc29, 32'hffd8dc29, 32'hffd8dc29, 32'hffd8dc29, 32'hff191919, 32'hff191919, 32'hffb002d7, 32'hffb002d7, 32'hff191919, 32'hff191919, 32'hffd8dc29, 32'hffd8dc29, 32'hffd8dc29, 32'hffd8dc29, 32'hff191919, 32'hffb002d7, 32'hff191919, 32'hff191919, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 
32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'hff191919, 32'hff191919, 32'hff191919, 32'hffd8dc29, 32'hffd8dc29, 32'hffd8dc29, 32'hffd8dc29, 32'hffd8dc29, 32'hff191919, 32'hffb002d7, 32'hffb002d7, 32'hff191919, 32'hffd8dc29, 32'hffd8dc29, 32'hffd8dc29, 32'hffd8dc29, 32'hffd8dc29, 32'hff191919, 32'hff191919, 32'hff191919, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 
32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'hff191919, 32'hff191919, 32'hff191919, 32'hffd8dc29, 32'hffd8dc29, 32'hffd8dc29, 32'hffd8dc29, 32'hff191919, 32'hff191919, 32'hff191919, 32'hff191919, 32'hffd8dc29, 32'hffd8dc29, 32'hffd8dc29, 32'hffd8dc29, 32'hff191919, 32'hff191919, 32'hff191919, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 
32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'hff191919, 32'hffd8dc29, 32'hffd8dc29, 32'hffd8dc29, 32'hffd8dc29, 32'hffd8dc29, 32'hff191919, 32'hff191919, 32'hffd8dc29, 32'hffd8dc29, 32'hffd8dc29, 32'hffd8dc29, 32'hffd8dc29, 32'hff191919, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 
32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'hff191919, 32'hffd8dc29, 32'hffd8dc29, 32'hffd8dc29, 32'hffd8dc29, 32'hffd8dc29, 32'hff191919, 32'hff191919, 32'hffd8dc29, 32'hffd8dc29, 32'hffd8dc29, 32'hffd8dc29, 32'hffd8dc29, 32'hff191919, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 
32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'hff191919, 32'hffd8dc29, 32'hff191919, 32'hff191919, 32'hff191919, 32'hffd8dc29, 32'hffd8dc29, 32'hffd8dc29, 32'hffd8dc29, 32'hff191919, 32'hff191919, 32'hff191919, 32'hff191919, 32'hff191919, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 
32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'hff191919, 32'hff191919, 32'hffffffff, 32'hffffffff, 32'hffffffff, 32'hff191919, 32'hffd8dc29, 32'hffd8dc29, 32'hff191919, 32'hffffffff, 32'hffffffff, 32'hffffffff, 32'hff191919, 32'hff191919, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 
32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'hff191919, 32'hff191919, 32'hffffffff, 32'hff191919, 32'hff191919, 32'hff191919, 32'hffd8dc29, 32'hffd8dc29, 32'hff191919, 32'hff191919, 32'hff191919, 32'hffffffff, 32'hff191919, 32'hff191919, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 
32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'hff191919, 32'hffffffff, 32'hffffffff, 32'hff191919, 32'hff191919, 32'hffd8dc29, 32'hffd8dc29, 32'hff191919, 32'hff191919, 32'hffffffff, 32'hffffffff, 32'hff191919, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 
32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'hff191919, 32'hff191919, 32'hff191919, 32'hff191919, 32'hff191919, 32'hffd8dc29, 32'hffd8dc29, 32'hffd8dc29, 32'hff191919, 32'hff191919, 32'hff191919, 32'hff191919, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 
32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'hff191919, 32'hffd8dc29, 32'hffd8dc29, 32'hffd8dc29, 32'hffd8dc29, 32'hffd8dc29, 32'hffd8dc29, 32'hffd8dc29, 32'hffd8dc29, 32'hff191919, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 
32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'hff191919, 32'hff191919, 32'hff191919, 32'hffd8dc29, 32'hffd8dc29, 32'hffd8dc29, 32'hffd8dc29, 32'hff191919, 32'hff191919, 32'hff191919, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 
32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'hff191919, 32'hff191919, 32'hff191919, 32'hff191919, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 
32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000
};
jodi_down = '{
32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 
32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'hff191919, 32'hff191919, 32'hff191919, 32'hff191919, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 
32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'hff191919, 32'hff191919, 32'hff191919, 32'hffd8dc29, 32'hffd8dc29, 32'hffd8dc29, 32'hffd8dc29, 32'hff191919, 32'hff191919, 32'hff191919, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 
32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'hff191919, 32'hffd8dc29, 32'hffd8dc29, 32'hffd8dc29, 32'hffd8dc29, 32'hffd8dc29, 32'hffd8dc29, 32'hffd8dc29, 32'hffd8dc29, 32'hff191919, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 
32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'hff191919, 32'hff191919, 32'hff191919, 32'hff191919, 32'hffd8dc29, 32'hffd8dc29, 32'hffd8dc29, 32'hff191919, 32'hff191919, 32'hff191919, 32'hff191919, 32'hff191919, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 
32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'hff191919, 32'hffffffff, 32'hffffffff, 32'hff191919, 32'hff191919, 32'hffd8dc29, 32'hffd8dc29, 32'hff191919, 32'hff191919, 32'hffffffff, 32'hffffffff, 32'hff191919, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 
32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'hff191919, 32'hff191919, 32'hffffffff, 32'hff191919, 32'hff191919, 32'hff191919, 32'hffd8dc29, 32'hffd8dc29, 32'hff191919, 32'hff191919, 32'hff191919, 32'hffffffff, 32'hff191919, 32'hff191919, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 
32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'hff191919, 32'hff191919, 32'hffffffff, 32'hffffffff, 32'hffffffff, 32'hff191919, 32'hffd8dc29, 32'hffd8dc29, 32'hff191919, 32'hffffffff, 32'hffffffff, 32'hffffffff, 32'hff191919, 32'hff191919, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 
32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'hff191919, 32'hff191919, 32'hff191919, 32'hff191919, 32'hff191919, 32'hffd8dc29, 32'hffd8dc29, 32'hffd8dc29, 32'hffd8dc29, 32'hff191919, 32'hff191919, 32'hff191919, 32'hffd8dc29, 32'hff191919, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 
32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'hff191919, 32'hffd8dc29, 32'hffd8dc29, 32'hffd8dc29, 32'hffd8dc29, 32'hffd8dc29, 32'hff191919, 32'hff191919, 32'hffd8dc29, 32'hffd8dc29, 32'hffd8dc29, 32'hffd8dc29, 32'hffd8dc29, 32'hff191919, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 
32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'hff191919, 32'hffd8dc29, 32'hffd8dc29, 32'hffd8dc29, 32'hffd8dc29, 32'hffd8dc29, 32'hff191919, 32'hff191919, 32'hffd8dc29, 32'hffd8dc29, 32'hffd8dc29, 32'hffd8dc29, 32'hffd8dc29, 32'hff191919, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 
32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'hff191919, 32'hff191919, 32'hff191919, 32'hffd8dc29, 32'hffd8dc29, 32'hffd8dc29, 32'hffd8dc29, 32'hff191919, 32'hff191919, 32'hff191919, 32'hff191919, 32'hffd8dc29, 32'hffd8dc29, 32'hffd8dc29, 32'hffd8dc29, 32'hff191919, 32'hff191919, 32'hff191919, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 
32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'hff191919, 32'hff191919, 32'hff191919, 32'hffd8dc29, 32'hffd8dc29, 32'hffd8dc29, 32'hffd8dc29, 32'hffd8dc29, 32'hff191919, 32'hffb002d7, 32'hffb002d7, 32'hff191919, 32'hffd8dc29, 32'hffd8dc29, 32'hffd8dc29, 32'hffd8dc29, 32'hffd8dc29, 32'hff191919, 32'hff191919, 32'hff191919, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 
32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'hff191919, 32'hff191919, 32'hffb002d7, 32'hff191919, 32'hffd8dc29, 32'hffd8dc29, 32'hffd8dc29, 32'hffd8dc29, 32'hff191919, 32'hff191919, 32'hffb002d7, 32'hffb002d7, 32'hff191919, 32'hff191919, 32'hffd8dc29, 32'hffd8dc29, 32'hffd8dc29, 32'hffd8dc29, 32'hff191919, 32'hffb002d7, 32'hff191919, 32'hff191919, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 
32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'hff191919, 32'hffb002d7, 32'hffb002d7, 32'hff191919, 32'hffd8dc29, 32'hffd8dc29, 32'hffd8dc29, 32'hffd8dc29, 32'hff191919, 32'hffb002d7, 32'hffb002d7, 32'hffb002d7, 32'hffb002d7, 32'hff191919, 32'hffd8dc29, 32'hffd8dc29, 32'hffd8dc29, 32'hffd8dc29, 32'hff191919, 32'hffb002d7, 32'hffb002d7, 32'hff191919, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 
32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'hff191919, 32'hffb002d7, 32'hffb002d7, 32'hff191919, 32'hffd8dc29, 32'hffd8dc29, 32'hffd8dc29, 32'hffd8dc29, 32'hff191919, 32'hffb002d7, 32'hffb002d7, 32'hffb002d7, 32'hffb002d7, 32'hff191919, 32'hffd8dc29, 32'hffd8dc29, 32'hffd8dc29, 32'hffd8dc29, 32'hff191919, 32'hffb002d7, 32'hffb002d7, 32'hff191919, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 
32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'hff191919, 32'hff191919, 32'hffb002d7, 32'hffb002d7, 32'hff191919, 32'hffd8dc29, 32'hffd8dc29, 32'hffd8dc29, 32'hffd8dc29, 32'hff191919, 32'hffb002d7, 32'hffb002d7, 32'hffb002d7, 32'hffb002d7, 32'hff191919, 32'hffd8dc29, 32'hffd8dc29, 32'hffd8dc29, 32'hffd8dc29, 32'hff191919, 32'hffb002d7, 32'hffb002d7, 32'hff191919, 32'hff191919, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 
32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'hff191919, 32'hffb002d7, 32'hffb002d7, 32'hffb002d7, 32'hff191919, 32'hffd8dc29, 32'hffd8dc29, 32'hffd8dc29, 32'hffd8dc29, 32'hff191919, 32'hffb002d7, 32'hffb002d7, 32'hffb002d7, 32'hffb002d7, 32'hff191919, 32'hffd8dc29, 32'hffd8dc29, 32'hffd8dc29, 32'hffd8dc29, 32'hff191919, 32'hffb002d7, 32'hffb002d7, 32'hffb002d7, 32'hff191919, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 
32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'hff191919, 32'hffb002d7, 32'hffb002d7, 32'hffb002d7, 32'hff191919, 32'hffd8dc29, 32'hffd8dc29, 32'hffd8dc29, 32'hffd8dc29, 32'hff191919, 32'hff191919, 32'hffb002d7, 32'hffb002d7, 32'hff191919, 32'hff191919, 32'hffd8dc29, 32'hffd8dc29, 32'hffd8dc29, 32'hffd8dc29, 32'hff191919, 32'hffb002d7, 32'hffb002d7, 32'hffb002d7, 32'hff191919, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 
32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'hff191919, 32'hff191919, 32'hff191919, 32'hffb002d7, 32'hff191919, 32'hffd8dc29, 32'hffd8dc29, 32'hffd8dc29, 32'hffd8dc29, 32'hffd8dc29, 32'hff191919, 32'hffb002d7, 32'hffb002d7, 32'hff191919, 32'hffd8dc29, 32'hffd8dc29, 32'hffd8dc29, 32'hffd8dc29, 32'hffd8dc29, 32'hff191919, 32'hffb002d7, 32'hff191919, 32'hff191919, 32'hff191919, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 
32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'hff191919, 32'hff191919, 32'hff191919, 32'hff191919, 32'hffd8dc29, 32'hffd8dc29, 32'hffd8dc29, 32'hffd8dc29, 32'hff191919, 32'hffb002d7, 32'hffb002d7, 32'hff191919, 32'hffd8dc29, 32'hffd8dc29, 32'hffd8dc29, 32'hffd8dc29, 32'hff191919, 32'hff191919, 32'hff191919, 32'hff191919, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 
32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'hff191919, 32'hff191919, 32'hffd8dc29, 32'hffd8dc29, 32'hffd8dc29, 32'hff191919, 32'hff191919, 32'hff191919, 32'hff191919, 32'hffd8dc29, 32'hffd8dc29, 32'hffd8dc29, 32'hff191919, 32'hff191919, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 
32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'hff191919, 32'hff191919, 32'hffd8dc29, 32'hffd8dc29, 32'hffd8dc29, 32'hff191919, 32'hff191919, 32'hffd8dc29, 32'hffd8dc29, 32'hffd8dc29, 32'hff191919, 32'hff191919, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 
32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'hff191919, 32'hff191919, 32'hffd8dc29, 32'hffd8dc29, 32'hffd8dc29, 32'hffd8dc29, 32'hffd8dc29, 32'hffd8dc29, 32'hff191919, 32'hff191919, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 
32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'hff191919, 32'hff191919, 32'hffd8dc29, 32'hffd8dc29, 32'hffd8dc29, 32'hffd8dc29, 32'hff191919, 32'hff191919, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 
32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'hff191919, 32'hff191919, 32'hffd8dc29, 32'hffd8dc29, 32'hff191919, 32'hff191919, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 
32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'hff191919, 32'hffd8dc29, 32'hffd8dc29, 32'hff191919, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 
32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'hff191919, 32'hff191919, 32'hff191919, 32'hffd8dc29, 32'hffd8dc29, 32'hff191919, 32'hff191919, 32'hff191919, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 
32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'hff191919, 32'hff191919, 32'hffd8dc29, 32'hffb002d7, 32'hffd8dc29, 32'hffb002d7, 32'hffd8dc29, 32'hffd8dc29, 32'hff191919, 32'hff191919, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 
32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'hff191919, 32'hff191919, 32'hffb002d7, 32'hffd8dc29, 32'hffb002d7, 32'hffb002d7, 32'hffd8dc29, 32'hffb002d7, 32'hffb002d7, 32'hffd8dc29, 32'hffb002d7, 32'hffb002d7, 32'hff191919, 32'hff191919, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 
32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'hff191919, 32'hff191919, 32'hffb002d7, 32'hffb002d7, 32'hffb002d7, 32'hffd8dc29, 32'hffb002d7, 32'hffb002d7, 32'hffd8dc29, 32'hffb002d7, 32'hffb002d7, 32'hffd8dc29, 32'hffd8dc29, 32'hffd8dc29, 32'hffb002d7, 32'hffb002d7, 32'hff191919, 32'hff191919, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 
32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'hff191919, 32'hff191919, 32'hff191919, 32'hff191919, 32'hff191919, 32'hff191919, 32'hff191919, 32'hff191919, 32'hff191919, 32'hff191919, 32'hff191919, 32'hff191919, 32'hff191919, 32'hff191919, 32'hff191919, 32'hff191919, 32'hff191919, 32'hff191919, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000
};

	Xval = X;
	Yval = Y;
end

always_ff @(posedge frame_clk)
begin
	color <= 32'h00000000;
	unique case(last_key_code)//unique-16 case(keycode[7:0])
	//jodi_left	
	8'h50: 
	begin
	color <= jodi_left [Yval*32+Xval];
	end
	//jodi_right
	8'h4F: 
	begin
	color <= jodi_right [Yval*32+Xval];
	end
	//jodi_up
	8'h52: 
	begin
	color <= jodi_up [Yval*32+Xval];
	end
	//jodi_down
	8'h51: 
	begin
	color <= jodi_down [Yval*32+Xval];
	end	
	default:;
	endcase
end


endmodule
